`timescale 1ns/1ns
module TM_Pipeline();

    reg clk, rst;

    initial begin
        clk = 1;
	forever #5 clk = ~clk;
    end

    initial begin
	rst = 1'b1;
	$readmemh("instr_mem.txt", CPU.instrMem.mem_array );
	$readmemh("data_mem.txt", CPU.dataMemory.mem_array );
	$readmemh("reg.txt", CPU.regFile.file_array );
	#10;
	rst = 1'b0;
    end
    always @( posedge clk ) begin
	
        $display( "%d, PC:", $time/10-1, CPU.pc );

	if ( CPU.op_code == 6'd0 ) begin

	    $display( "%d, wd: %d", $time/10-1, CPU.wb_wd );

	    if ( CPU.funct == 6'd32 ) $display( "%d, ADD\n", $time/10-1 );
	    else if ( CPU.funct == 6'd34 ) $display( "%d, SUB\n", $time/10-1 );
	    else if ( CPU.funct == 6'd36 ) $display( "%d, AND\n", $time/10-1 );
	    else if ( CPU.funct == 6'd37 ) $display( "%d, OR\n", $time/10-1 );
            else if ( CPU.funct == 6'd13 ) $display( "%d, ORI\n", $time/10-1 );
            else if ( CPU.funct == 6'd0 ) $display( "%d, NOP\n", $time/10-1 );
	end
        else if ( CPU.op_code == 6'd35 ) $display( "%d, LW\n", $time/10-1 );
        else if ( CPU.op_code == 6'd43 ) $display( "%d, SW\n", $time/10-1 );
	else if ( CPU.op_code == 6'd4 ) $display( "%d, BEQ\n", $time/10-1 );
	else if ( CPU.op_code == 6'd2 ) $display( "%d, J\n", $time/10-1 );
    end
	
    Pipeline_CPU CPU( clk, rst );
    
endmodule
